module wallace_tree(

);

endmodule
