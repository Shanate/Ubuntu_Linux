module test()

endmodule
